library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity sigGen is
	generic(  
           BITS : natural := 16
           );
	port(  
            pOut : out std_logic_vector(BITS-1 downto 0);
            pClk : in std_logic
        );
end entity sigGen;

architecture sinc of sigGen is
    type integer_array is array (natural range<>) of integer;
    constant sinc_16 : integer_array (0 to 255) := (10876,10681,10641,10766,11039,11422,11860,12288,12643,12870,12934,12821,12547,12148,11682,11218,10824,10561,10471,10569,10845,11261,11757,12262,12699,13003,13125,13043,12767,12332,11801,11251,10764,10413,10254,10315,10592,11047,11618,12220,12766,13172,13374,13337,13061,12582,11966,11302,10688,10217,9963,9970,10243,10749,11419,12156,12853,13403,13721,13751,13482,12944,12210,11384,10586,9937,9539,9460,9723,10299,11113,12051,12978,13753,14255,14397,14146,13523,12607,11523,10427,9484,8841,8609,8842,9525,10578,11860,13190,14370,15214,15578,15380,14617,13371,11801,10123,8583,7423,6843,6974,7846,9387,11418,13671,15828,17554,18547,18584,17559,15508,12619,9219,5750,2720,648,0,1132,4238,9317,16157,24349,33317,42371,50772,57813,62883,65535,65535,62883,57813,50772,42371,33317,24349,16157,9317,4238,1132,0,648,2720,5750,9219,12619,15508,17559,18584,18547,17554,15828,13671,11418,9387,7846,6974,6843,7423,8583,10123,11801,13371,14617,15380,15578,15214,14370,13190,11860,10578,9525,8842,8609,8841,9484,10427,11523,12607,13523,14146,14397,14255,13753,12978,12051,11113,10299,9723,9460,9539,9937,10586,11384,12210,12944,13482,13751,13721,13403,12853,12156,11419,10749,10243,9970,9963,10217,10688,11302,11966,12582,13061,13337,13374,13172,12766,12220,11618,11047,10592,10315,10254,10413,10764,11251,11801,12332,12767,13043,13125,13003,12699,12262,11757,11261,10845,10569,10471,10561,10824,11218,11682,12148,12547,12821,12934,12870,12643,12288,11860,11422,11039,10766,10641,10681,10876); 
    signal addr,addr_i : std_logic_vector(7 downto 0) := (others=>'0');
begin

    process (pClk)
    begin
        if rising_edge(pClk) then
            pOut <= std_logic_vector(to_unsigned(sinc_16(to_integer(unsigned(addr))),BITS));
            addr <= addr_i;
        end if;
    end process;

    addr_i <= std_logic_vector(unsigned(addr)+to_unsigned(1,addr'length));

end architecture sinc;





