

package constants is
    constant  COMMAND_OSC_FAIL : integer := 255;
    constant  COMMAND_OSC_START : integer := 1;
    constant  COMMAND_OSC_DATA : integer := 2;
    constant  COMMAND_OSC_TLEVEL : integer := 3;
    constant  COMMAND_OSC_TEDGE : integer := 4;
    constant  COMMAND_OSC_STATUS : integer := 5;
end package constants;





