

package constants is
    constant  COMMAND_FAIL : integer := 255;
    constant  COMMAND_OSC_START : integer := 1;
    constant  COMMAND_OSC_DATA : integer := 2;
    constant  COMMAND_OSC_TLEVEL : integer := 3;
    constant  COMMAND_OSC_TEDGE : integer := 4;
    constant  COMMAND_OSC_STATUS : integer := 5;
    
    constant  COMMAND_HIST_START : integer := 6;
    constant  COMMAND_HIST_STOP : integer := 7;
    constant  COMMAND_HIST_DATA : integer := 8;
    constant  COMMAND_HIST_CLEAR : integer := 9;
    constant  COMMAND_HIST_TIME : integer := 10;
    constant  COMMAND_HIST_STATUS : integer := 11;

end package constants;





